module semaforo(A, B, VERA, VERB, VERMA, VERMB);

    input A, B;
    output VERA, VERB, VERMA, VERMB;

    assign VERA = 
    assign VERB =
    assign VERMA =
    assign VERMB =

endmodule